���      �sklearn.linear_model._base��LinearRegression���)��}�(�fit_intercept���copy_X���n_jobs�N�positive���n_features_in_�K�coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�C�Bs8S~?&#JN�D�?�t�b�rank_�K�	singular_�hhK ��h��R�(KK��h�C¨����U@�RtVU@�t�b�
intercept_�h�scalar���hC�v�����?���R��_sklearn_version��1.3.0�ub.